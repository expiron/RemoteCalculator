module RemoteCalculator(
	input            clk,
	input            reset,
	input      [3:0] row,
	input            rxd,
	output     [3:0] col,
	output     [3:0] com,
	output     [7:0] seg,
	output           txd,
	output           sign,
	output           clcZero
);

endmodule